Vim�UnDo� ��Oow�x~CF�.���ơJB���   s   module test_top();                             Yg�y    _�                             ����                                                                                                                                                                                                                                                                                                                                                             Yg�x    �         s      module test_top();5��