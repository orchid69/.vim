Vim�UnDo� |�O�יC��;2��sm`�o1��0O�   �           
      V       V   V   V    Y[�T    _�                             ����                                                                                                                                                                                                                                                                                                                                                             Y[��    �          �      module adjust_v(/*AUTOARG*/5�_�      !              �        ����                                                                                                                                                                                                                                                                                                                            �           �          v       Y[�w    �   �   �          	end�   �   �          		else s2_v_reg <= s1_v_reg;�   �   �          		if (!xrst) s2_v_reg <= 8'b0;�   �   �          ,	always @(posedge clk or negedge xrst) begin�   �   �           �   �   �          	end�   �   �          &		else s2_from_v_reg <= s1_from_v_reg;�   �   �          #		if (!xrst) s2_from_v_reg <= 8'b0;�   �   �          ,	always @(posedge clk or negedge xrst) begin�   �   �           �   �   �          	end�   �   �           		else s2_ack_reg <= s1_ack_reg;�   �   �           		if (!xrst) s2_ack_reg <= 1'b0;�   �   �          ,	always @(posedge clk or negedge xrst) begin�   �   �           �   �   �          	end�   �   �          *		else s2_quotient_s_reg <= s2_quotient_s;�   �   �          '		if (!xrst) s2_quotient_s_reg <= 8'd0;�   �   �          ,	always @(posedge clk or negedge xrst) begin�   �   �           �   �   �          	end�   �   �          *		else s2_quotient_l_reg <= s2_quotient_l;�   �   �          '		if (!xrst) s2_quotient_l_reg <= 8'd0;�   �   �          ,	always @(posedge clk or negedge xrst) begin5�_�       "           !   v       ����                                                                                                                                                                                                                                                                                                                            v          v          V       Y[�~     �   u   w          	reg [7:0] s2_quotient_l_reg;5�_�   !   #           "   w       ����                                                                                                                                                                                                                                                                                                                            w          w          V       Y[�    �   v   x          	reg [7:0] s2_quotient_s_reg;5�_�   "   $           #   u       ����                                                                                                                                                                                                                                                                                                                            u          u          V       Y[��     �   t   v          	reg s2_ack_reg;5�_�   #   %           $   y       ����                                                                                                                                                                                                                                                                                                                            y          y          V       Y[��     �   x   z          	reg [7:0] s2_from_v_reg;5�_�   $   &           %   z       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   y   {          	reg [7:0] s2_v_reg;5�_�   %   '           &   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      	reg [7:0] 	s3_v_reg;5�_�   &   (           '   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      	reg 		s3_ack_reg;5�_�   '   )           (   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      #	wire [7:0]      s3_quotient_l_sel;5�_�   (   *           )   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      #	wire [7:0]      s3_quotient_s_sel;5�_�   )   +           *   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      !	wire [7:0]      s3_quotient_sel;5�_�   *   ,           +   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      	wire [7:0]      s3_v;5�_�   +   -           ,   �   	    ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      O	assign s3_quotient_s_sel = (s2_from_v_reg != 8'd0) ? s2_quotient_s_reg : 8'd0;5�_�   ,   .           -   �   	    ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      Q	assign s3_quotient_l_sel = (s2_from_v_reg != 8'd255) ? s2_quotient_l_reg : 8'd0;5�_�   -   /           .   �   	    ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      ]	assign s3_quotient_sel = (s2_v_reg > s2_from_v_reg) ? s3_quotient_l_sel : s3_quotient_s_sel;5�_�   .   0           /   �   	    ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      E	assign s3_v = (s3_quotient_sel > 8'd255) ? 8'd255 : s3_quotient_sel;5�_�   /   1           0   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[�5     �   �   �   �      O	assign s2_quotient_s_sel = (s2_from_v_reg != 8'd0) ? s2_quotient_s_reg : 8'd0;5�_�   0   2           1   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[�5     �   �   �   �      Q	assign s2_quotient_l_sel = (s2_from_v_reg != 8'd255) ? s2_quotient_l_reg : 8'd0;5�_�   1   3           2   �   '    ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[�=     �   �   �   �      ]	assign s2_quotient_sel = (s2_v_reg > s2_from_v_reg) ? s3_quotient_l_sel : s3_quotient_s_sel;5�_�   2   4           3   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[�^     �   �   �   �      ]	assign s2_quotient_sel = (s2_v_reg > s1_from_v_reg) ? s3_quotient_l_sel : s3_quotient_s_sel;5�_�   3   5           4   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[�j     �   �   �   �      E	assign s2_v = (s3_quotient_sel > 8'd255) ? 8'd255 : s3_quotient_sel;5�_�   4   6           5   �   G    ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[�     �   �   �   �      O	assign s2_quotient_s_sel = (s1_from_v_reg != 8'd0) ? s2_quotient_s_reg : 8'd0;5�_�   5   7           6   �   I    ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[�     �   �   �   �      Q	assign s2_quotient_l_sel = (s1_from_v_reg != 8'd255) ? s2_quotient_l_reg : 8'd0;5�_�   6   8           7   �   8    ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[�     �   �   �   �      ]	assign s2_quotient_sel = (s1_v_reg > s1_from_v_reg) ? s3_quotient_l_sel : s3_quotient_s_sel;5�_�   7   9           8   �   L    ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      ]	assign s2_quotient_sel = (s1_v_reg > s1_from_v_reg) ? s2_quotient_l_sel : s3_quotient_s_sel;5�_�   8   :           9   �   6    ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      E	assign s2_v = (s2_quotient_sel > 8'd255) ? 8'd255 : s3_quotient_sel;5�_�   9   ;           :   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      		if (!xrst) s3_v_reg <= 8'd0;5�_�   :   <           ;   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      		else s3_v_reg <= s3_v;5�_�   ;   =           <   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      		else s2_v_reg <= s3_v;5�_�   <   >           =   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �       		if (!xrst) s3_ack_reg <= 1'b0;5�_�   =   ?           >   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �       		else s3_ack_reg <= s2_ack_reg;5�_�   >   @           ?   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��     �   �   �   �      	assign pixel_v_out = s3_v_reg;5�_�   ?   A           @   �       ����                                                                                                                                                                                                                                                                                                                            z          z          V       Y[��    �   �   �   �      	assign snd_ack = s3_ack_reg;5�_�   @   B           A   |       ����                                                                                                                                                                                                                                                                                                                                                             Y[��     �   {   }   �      	wire [7:0] s2_quotient_l;5�_�   A   C           B   }       ����                                                                                                                                                                                                                                                                                                                                                             Y[��     �   |   ~   �      	wire [7:0] s2_quotient_s;5�_�   B   D           C   �       ����                                                                                                                                                                                                                                                                                                                                                             Y[��     �   �   �   �      +			      .o1		(s2_quotient_l), // Templated5�_�   C   E           D   �       ����                                                                                                                                                                                                                                                                                                                                                             Y[�     �   �   �   �      +			      .o1		(s2_quotient_s), // Templated5�_�   D   F           E   �   7    ����                                                                                                                                                                                                                                                                                                                                                             Y[�     �   �   �   �      K	assign s2_quotient_s_sel = (s1_from_v_reg != 8'd0) ? s2_quotient_s : 8'd0;5�_�   E   G           F   �   9    ����                                                                                                                                                                                                                                                                                                                                                             Y[�   	 �   �   �   �      M	assign s2_quotient_l_sel = (s1_from_v_reg != 8'd255) ? s2_quotient_l : 8'd0;5�_�   F   H           G   �       ����                                                                                                                                                                                                                                                                                                                                                             Y[�     �   �   �   �       		else s2_ack_reg <= s2_ack_reg;5�_�   G   I           H   �   
    ����                                                                                                                                                                                                                                                                                                                                                             Y[�)     �   �   �   �      	// stage 3 (calculation3)5�_�   H   J           I   �       ����                                                                                                                                                                                                                                                                                                                                                             Y[�,     �   �   �   �      	// stage 2 (calculation3)5�_�   I   K           J   �        ����                                                                                                                                                                                                                                                                                                                            �           �           V        Y[�3     �   �   �          /	// always @(posedge clk or negedge xrst) begin   *	// 	if (!xrst) s2_quotient_l_reg <= 8'd0;   -	// 	else s2_quotient_l_reg <= s2_quotient_l;   	// end       //   /	// always @(posedge clk or negedge xrst) begin   *	// 	if (!xrst) s2_quotient_s_reg <= 8'd0;   -	// 	else s2_quotient_s_reg <= s2_quotient_s;   	// end       //   /	// always @(posedge clk or negedge xrst) begin   #	// 	if (!xrst) s2_ack_reg <= 1'b0;   #	// 	else s2_ack_reg <= s1_ack_reg;   	// end       //   /	// always @(posedge clk or negedge xrst) begin   &	// 	if (!xrst) s2_from_v_reg <= 8'b0;   )	// 	else s2_from_v_reg <= s1_from_v_reg;   	// end       //   /	// always @(posedge clk or negedge xrst) begin   !	// 	if (!xrst) s2_v_reg <= 8'b0;   	// 	else s2_v_reg <= s1_v_reg;   	// end    5�_�   J   L           K   r        ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�?     �   q   r          ;	//////////////////////////////////////////////////////////5�_�   K   M           L   r       ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�?     �   q   r          	// stage 2 (calculation2)5�_�   L   N           M   r       ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�?     �   q   r          ;	//////////////////////////////////////////////////////////5�_�   M   O           N   r       ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�?     �   q   r          	// reg s2_ack_reg;5�_�   N   P           O   r       ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�?     �   q   r           	// reg [7:0] s2_quotient_l_reg;5�_�   O   Q           P   r       ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�@     �   q   r           	// reg [7:0] s2_quotient_s_reg;5�_�   P   R           Q   r        ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�B     �   q   r           5�_�   Q   S           R   r       ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�C     �   q   r          	// reg [7:0] s2_from_v_reg;5�_�   R   T           S   r       ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�D     �   q   r          	// reg [7:0] s2_v_reg;5�_�   S   U           T   r        ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�E     �   q   r           5�_�   T   V           U   �       ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�O     �   �   �          ;	//////////////////////////////////////////////////////////   	// stage 2 (calculation2)   ;	//////////////////////////////////////////////////////////5�_�   U               V   q        ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[�S    �   q   u   �    �   q   r   �    5�_�                   u       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[�U    �   t   v          	// reg s2_ack_reg;�   u   w           	// reg [7:0] s2_quotient_l_reg;�   v   x           	// reg [7:0] s2_quotient_s_reg;�   w   y              //�   x   z          	// reg [7:0] s2_from_v_reg;�   y   {          	// reg [7:0] s2_v_reg;�   z   |              //�   {   }          	// wire [7:0] s2_quotient_l;�   |   ~          	// wire [7:0] s2_quotient_s;�   }                 //�   ~   �          	// /* div_u AUTO_TEMPLATE (�      �          	//  .i1(s1_dividend_l_reg),�   �   �          	//  .i2(s1_divisor_l_reg),�   �   �          	//  .o1(s2_quotient_l),�   �   �          	// );*/�   �   �          &	// div_u #(16,8,8) div0 (/*AUTOINST*/�   �   �          	// 		      // Outputs�   �   �          .	// 		      .o1		(s2_quotient_l), // Templated�   �   �          	// 		      // Inputs�   �   �          2	// 		      .i1		(s1_dividend_l_reg), // Templated�   �   �          2	// 		      .i2		(s1_divisor_l_reg)); // Templated�   �   �              //�   �   �          	// /* div_u AUTO_TEMPLATE (�   �   �          	//  .i1(s1_dividend_s_reg),�   �   �          	//  .i2(s1_divisor_s_reg),�   �   �          	//  .o1(s2_quotient_s),�   �   �          	// );*/�   �   �          &	// div_u #(16,8,8) div1 (/*AUTOINST*/�   �   �          	// 		      // Outputs�   �   �          .	// 		      .o1		(s2_quotient_s), // Templated�   �   �          	// 		      // Inputs�   �   �          2	// 		      .i1		(s1_dividend_s_reg), // Templated�   �   �          2	// 		      .i2		(s1_divisor_s_reg)); // Templated�   �   �              //�   �   �          /	// always @(posedge clk or negedge xrst) begin�   �   �          *	// 	if (!xrst) s2_quotient_l_reg <= 8'd0;�   �   �          -	// 	else s2_quotient_l_reg <= s2_quotient_l;�   �   �          	// end�   �   �              //�   �   �          /	// always @(posedge clk or negedge xrst) begin�   �   �          *	// 	if (!xrst) s2_quotient_s_reg <= 8'd0;�   �   �          -	// 	else s2_quotient_s_reg <= s2_quotient_s;�   �   �          	// end�   �   �              //�   �   �          /	// always @(posedge clk or negedge xrst) begin�   �   �          #	// 	if (!xrst) s2_ack_reg <= 1'b0;�   �   �          #	// 	else s2_ack_reg <= s1_ack_reg;�   �   �          	// end�   �   �              //�   �   �          /	// always @(posedge clk or negedge xrst) begin�   �   �          &	// 	if (!xrst) s2_from_v_reg <= 8'b0;�   �   �          )	// 	else s2_from_v_reg <= s1_from_v_reg;�   �   �          	// end�   �   �              //�   �   �          /	// always @(posedge clk or negedge xrst) begin�   �   �          !	// 	if (!xrst) s2_v_reg <= 8'b0;�   �   �          	// 	else s2_v_reg <= s1_v_reg;�   �   �          	// end5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[�}     �   �   �   �      	reg [7:0] 	s2_v_reg;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[�     �   �   �   �      	reg 		s2_ack_reg;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ހ     �   �   �   �      #	wire [7:0]      s2_quotient_l_sel;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ށ     �   �   �   �      #	wire [7:0]      s2_quotient_s_sel;5�_�      	              �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ށ     �   �   �   �      !	wire [7:0]      s2_quotient_sel;5�_�      
           	   �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ނ     �   �   �   �      	wire [7:0]      s2_v;5�_�   	              
   �   	    ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ކ     �   �   �   �      O	assign s2_quotient_s_sel = (s2_from_v_reg != 8'd0) ? s2_quotient_s_reg : 8'd0;5�_�   
                 �   	    ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ކ     �   �   �   �      Q	assign s2_quotient_l_sel = (s2_from_v_reg != 8'd255) ? s2_quotient_l_reg : 8'd0;5�_�                    �   	    ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[އ     �   �   �   �      ]	assign s2_quotient_sel = (s2_v_reg > s2_from_v_reg) ? s3_quotient_l_sel : s3_quotient_s_sel;5�_�                    �   	    ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[އ     �   �   �   �      E	assign s2_v = (s3_quotient_sel > 8'd255) ? 8'd255 : s3_quotient_sel;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ދ     �   �   �   �      O	assign s2_quotient_s_sel = (s1_from_v_reg != 8'd0) ? s2_quotient_s_reg : 8'd0;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ތ     �   �   �   �      Q	assign s2_quotient_l_sel = (s1_from_v_reg != 8'd255) ? s2_quotient_l_reg : 8'd0;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ލ     �   �   �   �      ]	assign s2_quotient_sel = (s1_v_reg > s2_from_v_reg) ? s3_quotient_l_sel : s3_quotient_s_sel;5�_�                    �   '    ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ސ     �   �   �   �      ]	assign s2_quotient_sel = (s1_v_reg > s1_from_v_reg) ? s3_quotient_l_sel : s3_quotient_s_sel;5�_�                    �   7    ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ޓ     �   �   �   �      O	assign s2_quotient_s_sel = (s1_from_v_reg != 8'd0) ? s1_quotient_s_reg : 8'd0;5�_�                    �   9    ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ޔ     �   �   �   �      Q	assign s2_quotient_l_sel = (s1_from_v_reg != 8'd255) ? s1_quotient_l_reg : 8'd0;5�_�                    �   8    ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ަ     �   �   �   �      ]	assign s2_quotient_sel = (s1_v_reg > s1_from_v_reg) ? s2_quotient_l_sel : s3_quotient_s_sel;5�_�                    �   6    ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ާ     �   �   �   �      E	assign s2_v = (s3_quotient_sel > 8'd255) ? 8'd255 : s2_quotient_sel;5�_�                    �   L    ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[ު     �   �   �   �      ]	assign s2_quotient_sel = (s1_v_reg > s1_from_v_reg) ? s2_quotient_l_sel : s2_quotient_s_sel;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[޵     �   �   �   �      		if (!xrst) s2_v_reg <= 8'd0;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[޷     �   �   �   �       		if (!xrst) s2_ack_reg <= 1'b0;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[޼     �   �   �   �       		else s2_ack_reg <= s2_ack_reg;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[��     �   �   �   �       		else s2_ack_reg <= s1_ack_reg;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[��     �   �   �   �      E	assign s2_v = (s2_quotient_sel > 8'd255) ? 8'd255 : s2_quotient_sel;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[��     �   �   �   �      		else s2_v_reg <= s3_v;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[��     �   �   �   �      		else s2_v_reg <= s2_v;5�_�                    �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[��     �   �   �   �      	assign pixel_v_out = s2_v_reg;5�_�                     �       ����                                                                                                                                                                                                                                                                                                                            u          �          v       Y[��    �   �   �   �      	assign snd_ack = s2_ack_reg;5�_�                    �        ����                                                                                                                                                                                                                                                                                                                            �          �           V        Y[��     �   �   �          >	// //////////////////////////////////////////////////////////�   �   �          	// // stage 3 (calculation3)�   �   �          >	// //////////////////////////////////////////////////////////�   �   �          	// reg [7:0] 	s3_v_reg;�   �   �          	// reg 		s3_ack_reg;�   �   �          &	// wire [7:0]      s3_quotient_l_sel;�   �   �          &	// wire [7:0]      s3_quotient_s_sel;�   �   �          $	// wire [7:0]      s3_quotient_sel;�   �   �              //�   �   �          	// wire [7:0]      s3_v;�   �   �              //�   �   �          R	// assign s3_quotient_s_sel = (s2_from_v_reg != 8'd0) ? s2_quotient_s_reg : 8'd0;�   �   �          T	// assign s3_quotient_l_sel = (s2_from_v_reg != 8'd255) ? s2_quotient_l_reg : 8'd0;�   �   �          `	// assign s3_quotient_sel = (s2_v_reg > s2_from_v_reg) ? s3_quotient_l_sel : s3_quotient_s_sel;�   �   �          H	// assign s3_v = (s3_quotient_sel > 8'd255) ? 8'd255 : s3_quotient_sel;�   �   �              //�   �   �          /	// always @(posedge clk or negedge xrst) begin�   �   �          !	// 	if (!xrst) s3_v_reg <= 8'd0;�   �   �          	// 	else s3_v_reg <= s3_v;�   �   �          	// end�   �   �              //�   �   �          /	// always @(posedge clk or negedge xrst) begin�   �   �          #	// 	if (!xrst) s3_ack_reg <= 1'b0;�   �   �          #	// 	else s3_ack_reg <= s2_ack_reg;�   �   �          	// end�   �   �              //5��