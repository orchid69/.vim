Vim�UnDo� 2��UkG:�-<��6���;��3��!:�Sp�ca   G   module top(      
                       Y[ؐ    _�                         
    ����                                                                                                                                                                                                                                                                                                                                                             Y[؏    �          G      module top(5��