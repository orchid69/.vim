Vim�UnDo� �,ET�����C�����*����똮 �B=A��   G      adjust_v_2 adj0(// Outputs   /                          Y\�    _�                            ����                                                                                                                                                                                                                                                                                                                                                             Y\�    �          G      module top_2(5�_�                     /       ����                                                                                                                                                                                                                                                                                                                                                             Y\�    �   .   0   G         adjust_v_2 adj0(// Outputs5��