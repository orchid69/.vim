Vim�UnDo� pK����Jg�u�b�����k��P��@_{+�_K$   �   module adjust_v_2(/*AUTOARG*/                             Y[�1    _�                             ����                                                                                                                                                                                                                                                                                                                                                             Y[�0    �          �      module adjust_v_2(/*AUTOARG*/5��