Vim�UnDo� =--i�mS�����r���-ʄ���<~v   �      top_2 top0(// Outputs   V                          Y\j    _�                            ����                                                                                                                                                                                                                                                                                                                                                             Y\    �         �      module test_top_2();5�_�                    V       ����                                                                                                                                                                                                                                                                                                                                                             Y\i    �   U   W   �         top_2 top0(// Outputs5�_�                    V       ����                                                                                                                                                                                                                                                                                                                                                             Y\_     �   U   W   �         top_2 top0(// Outputs5��