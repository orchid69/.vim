Vim�UnDo� ���y���F�<� �k�Y-�8�d���gɧ6   �   module test_top();                             Y[إ    _�                             ����                                                                                                                                                                                                                                                                                                                                                             Y[ؤ    �         �      module test_top();5��